interface intf();
  logic d;
  logic q;
  logic qbar;
  logic clk;
  logic rst;
endinterface